// the below program is the and gate in the behavioral modeling
module andgate(
    input a,
    input b,
    output y
    );
    assign y = a&b;
endmodule
